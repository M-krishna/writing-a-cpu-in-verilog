module lc(
    
);
endmodule
