module my_basic_cpu;
    initial begin
	$display("Hello World");
    end
endmodule
