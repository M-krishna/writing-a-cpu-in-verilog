module my_basic_cpu_tb;
    my_basic_cpu mbc ();

    initial begin
	#5;
    end
endmodule
