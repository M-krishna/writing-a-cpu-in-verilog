module example;
    initial begin
	$display("Hello world");
    end
endmodule
