module example_tb;
    example e ();

    initial begin
	#1;
    end
endmodule
